library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity rom is
--  Port ( );
end rom;

architecture Behavioral of rom is

begin


end Behavioral;
