LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FSM IS
    --  Port ( );
    PORT (
        clk : IN STD_ULOGIC;
        VGA_DAddr : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
        data : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END FSM;